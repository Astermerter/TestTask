module main(
        input [15:0] first_num, // ��� �++ ������ ��������
        input [15:0] second_num, // ��� ����
        output reg [31:0] solution // � ���
);
        reg [3:0] n = 1; // ��� ������ ��� ���� ��������� �������
        reg [3:0] m;
        reg [15:0] F_F_P; // ������ ����� ������� �����
        reg [15:0] F_S_P; // ������ ����� ������� �����
        reg [15:0] S_F_P; // ���������� ������ �����
        reg [15:0] S_S_P;

        reg [15:0] p1;
        reg [15:0] p2;
        reg [15:0] p3;
        reg [15:0] p4;

        integer buf1; // (10^m) buf ���������������� ��� ��������� ����������
        integer buf2; // (10^2m)
        integer i;
        always @(*) begin
                if (n > 1) begin
                        m = n >> 1;
                        solution = 0;
                        buf1 = 10;
                        buf2 = 10;
                        for (i = 0; i < m - 1; i++) begin
                                buf1 = buf1 * 10;
                        end
                        for (i = 0; i < 2 * m - 1; i++) begin
                                buf2 = buf2 * 10;
                        end
                        F_F_P = first_num / buf1;
                        F_S_P = first_num % buf1;
                        S_F_P = second_num / buf1;
                        S_S_P = second_num % buf1;

                        p1 = F_F_P * S_F_P;
                        p2 = F_S_P * S_S_P;
                        p3 = (F_F_P + F_S_P)*(S_F_P + S_S_P);
                        p4 = p3 - p2 - p1;

                        solution = p1 * buf2 + p4 * buf1 + p2;
                end else begin
                        solution = first_num * second_num;
                end
        end
endmodule